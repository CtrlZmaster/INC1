library IEEE;
use IEEE.std_logic_1164.all;

package testbench_pkg is
   constant FILE_NAME : string := "chk_sim_sig_advanced.txt";

   constant N_TEST_WORDS : integer := 1676; 
   type t_test_words     is array (1 to N_TEST_WORDS) 
                                  of string(1 to 15);
   constant test_words : t_test_words :=
   ( 
     "0700146915#    ",
     "1700146915#    ",
     "2700146915#    ",
     "3700146915#    ",
     "4700146915#    ",
     "5700146915#    ",
     "6700146915#    ",
     "7700146915#    ",
     "8700146915#    ",
     "9700146915#    ",
     "A700146915#    ",
     "B700146915#    ",
     "C700146915#    ",
     "D700146915#    ",
     "*700146915#    ",
     "1000146915#    ",
     "1100146915#    ",
     "1200146915#    ",
     "1300146915#    ",
     "1400146915#    ",
     "1500146915#    ",
     "1600146915#    ",
     "1700146915#    ",
     "1800146915#    ",
     "1900146915#    ",
     "1A00146915#    ",
     "1B00146915#    ",
     "1C00146915#    ",
     "1D00146915#    ",
     "1*00146915#    ",
     "1700146915#    ",
     "1710146915#    ",
     "1720146915#    ",
     "1730146915#    ",
     "1740146915#    ",
     "1750146915#    ",
     "1760146915#    ",
     "1770146915#    ",
     "1780146915#    ",
     "1790146915#    ",
     "17A0146915#    ",
     "17B0146915#    ",
     "17C0146915#    ",
     "17D0146915#    ",
     "17*0146915#    ",
     "1700146915#    ",
     "1701146915#    ",
     "1702146915#    ",
     "1703146915#    ",
     "1704146915#    ",
     "1705146915#    ",
     "1706146915#    ",
     "1707146915#    ",
     "1708146915#    ",
     "1709146915#    ",
     "170A146915#    ",
     "170B146915#    ",
     "170C146915#    ",
     "170D146915#    ",
     "170*146915#    ",
     "1700046915#    ",
     "1700146915#    ",
     "1700246915#    ",
     "1700346915#    ",
     "1700446915#    ",
     "1700546915#    ",
     "1700646915#    ",
     "1700746915#    ",
     "1700846915#    ",
     "1700946915#    ",
     "1700A46915#    ",
     "1700B46915#    ",
     "1700C46915#    ",
     "1700D46915#    ",
     "1700*46915#    ",
     "1700106915#    ",
     "1700116915#    ",
     "1700126915#    ",
     "1700136915#    ",
     "1700146915#    ",
     "1700156915#    ",
     "1700166915#    ",
     "1700176915#    ",
     "1700186915#    ",
     "1700196915#    ",
     "17001A6915#    ",
     "17001B6915#    ",
     "17001C6915#    ",
     "17001D6915#    ",
     "17001*6915#    ",
     "1700140915#    ",
     "1700141915#    ",
     "1700142915#    ",
     "1700143915#    ",
     "1700144915#    ",
     "1700145915#    ",
     "1700146915#    ",
     "1700147915#    ",
     "1700148915#    ",
     "1700149915#    ",
     "170014A915#    ",
     "170014B915#    ",
     "170014C915#    ",
     "170014D915#    ",
     "170014*915#    ",
     "1700146015#    ",
     "1700146115#    ",
     "1700146215#    ",
     "1700146315#    ",
     "1700146415#    ",
     "1700146515#    ",
     "1700146615#    ",
     "1700146715#    ",
     "1700146815#    ",
     "1700146915#    ",
     "1700146A15#    ",
     "1700146B15#    ",
     "1700146C15#    ",
     "1700146D15#    ",
     "1700146*15#    ",
     "1700146905#    ",
     "1700146915#    ",
     "1700146925#    ",
     "1700146935#    ",
     "1700146945#    ",
     "1700146955#    ",
     "1700146965#    ",
     "1700146975#    ",
     "1700146985#    ",
     "1700146995#    ",
     "17001469A5#    ",
     "17001469B5#    ",
     "17001469C5#    ",
     "17001469D5#    ",
     "17001469*5#    ",
     "1700146910#    ",
     "1700146911#    ",
     "1700146912#    ",
     "1700146913#    ",
     "1700146914#    ",
     "1700146915#    ",
     "1700146916#    ",
     "1700146917#    ",
     "1700146918#    ",
     "1700146919#    ",
     "170014691A#    ",
     "170014691B#    ",
     "170014691C#    ",
     "170014691D#    ",
     "170014691*#    ",
     "00#            ",
     "01#            ",
     "02#            ",
     "03#            ",
     "04#            ",
     "05#            ",
     "06#            ",
     "07#            ",
     "08#            ",
     "09#            ",
     "0A#            ",
     "0B#            ",
     "0C#            ",
     "0D#            ",
     "0*#            ",
     "0#             ",
     "10#            ",
     "11#            ",
     "12#            ",
     "13#            ",
     "14#            ",
     "15#            ",
     "16#            ",
     "17#            ",
     "18#            ",
     "19#            ",
     "1A#            ",
     "1B#            ",
     "1C#            ",
     "1D#            ",
     "1*#            ",
     "1#             ",
     "20#            ",
     "21#            ",
     "22#            ",
     "23#            ",
     "24#            ",
     "25#            ",
     "26#            ",
     "27#            ",
     "28#            ",
     "29#            ",
     "2A#            ",
     "2B#            ",
     "2C#            ",
     "2D#            ",
     "2*#            ",
     "2#             ",
     "30#            ",
     "31#            ",
     "32#            ",
     "33#            ",
     "34#            ",
     "35#            ",
     "36#            ",
     "37#            ",
     "38#            ",
     "39#            ",
     "3A#            ",
     "3B#            ",
     "3C#            ",
     "3D#            ",
     "3*#            ",
     "3#             ",
     "40#            ",
     "41#            ",
     "42#            ",
     "43#            ",
     "44#            ",
     "45#            ",
     "46#            ",
     "47#            ",
     "48#            ",
     "49#            ",
     "4A#            ",
     "4B#            ",
     "4C#            ",
     "4D#            ",
     "4*#            ",
     "4#             ",
     "50#            ",
     "51#            ",
     "52#            ",
     "53#            ",
     "54#            ",
     "55#            ",
     "56#            ",
     "57#            ",
     "58#            ",
     "59#            ",
     "5A#            ",
     "5B#            ",
     "5C#            ",
     "5D#            ",
     "5*#            ",
     "5#             ",
     "60#            ",
     "61#            ",
     "62#            ",
     "63#            ",
     "64#            ",
     "65#            ",
     "66#            ",
     "67#            ",
     "68#            ",
     "69#            ",
     "6A#            ",
     "6B#            ",
     "6C#            ",
     "6D#            ",
     "6*#            ",
     "6#             ",
     "70#            ",
     "71#            ",
     "72#            ",
     "73#            ",
     "74#            ",
     "75#            ",
     "76#            ",
     "77#            ",
     "78#            ",
     "79#            ",
     "7A#            ",
     "7B#            ",
     "7C#            ",
     "7D#            ",
     "7*#            ",
     "7#             ",
     "80#            ",
     "81#            ",
     "82#            ",
     "83#            ",
     "84#            ",
     "85#            ",
     "86#            ",
     "87#            ",
     "88#            ",
     "89#            ",
     "8A#            ",
     "8B#            ",
     "8C#            ",
     "8D#            ",
     "8*#            ",
     "8#             ",
     "90#            ",
     "91#            ",
     "92#            ",
     "93#            ",
     "94#            ",
     "95#            ",
     "96#            ",
     "97#            ",
     "98#            ",
     "99#            ",
     "9A#            ",
     "9B#            ",
     "9C#            ",
     "9D#            ",
     "9*#            ",
     "9#             ",
     "A0#            ",
     "A1#            ",
     "A2#            ",
     "A3#            ",
     "A4#            ",
     "A5#            ",
     "A6#            ",
     "A7#            ",
     "A8#            ",
     "A9#            ",
     "AA#            ",
     "AB#            ",
     "AC#            ",
     "AD#            ",
     "A*#            ",
     "A#             ",
     "B0#            ",
     "B1#            ",
     "B2#            ",
     "B3#            ",
     "B4#            ",
     "B5#            ",
     "B6#            ",
     "B7#            ",
     "B8#            ",
     "B9#            ",
     "BA#            ",
     "BB#            ",
     "BC#            ",
     "BD#            ",
     "B*#            ",
     "B#             ",
     "C0#            ",
     "C1#            ",
     "C2#            ",
     "C3#            ",
     "C4#            ",
     "C5#            ",
     "C6#            ",
     "C7#            ",
     "C8#            ",
     "C9#            ",
     "CA#            ",
     "CB#            ",
     "CC#            ",
     "CD#            ",
     "C*#            ",
     "C#             ",
     "D0#            ",
     "D1#            ",
     "D2#            ",
     "D3#            ",
     "D4#            ",
     "D5#            ",
     "D6#            ",
     "D7#            ",
     "D8#            ",
     "D9#            ",
     "DA#            ",
     "DB#            ",
     "DC#            ",
     "DD#            ",
     "D*#            ",
     "D#             ",
     "*0#            ",
     "*1#            ",
     "*2#            ",
     "*3#            ",
     "*4#            ",
     "*5#            ",
     "*6#            ",
     "*7#            ",
     "*8#            ",
     "*9#            ",
     "*A#            ",
     "*B#            ",
     "*C#            ",
     "*D#            ",
     "**#            ",
     "*#             ",
     "1700146900#    ",
     "1700146901#    ",
     "1700146902#    ",
     "1700146903#    ",
     "1700146904#    ",
     "1700146905#    ",
     "1700146906#    ",
     "1700146907#    ",
     "1700146908#    ",
     "1700146909#    ",
     "170014690A#    ",
     "170014690B#    ",
     "170014690C#    ",
     "170014690D#    ",
     "170014690*#    ",
     "170014690#     ",
     "1700146910#    ",
     "1700146911#    ",
     "1700146912#    ",
     "1700146913#    ",
     "1700146914#    ",
     "1700146915#    ",
     "1700146916#    ",
     "1700146917#    ",
     "1700146918#    ",
     "1700146919#    ",
     "170014691A#    ",
     "170014691B#    ",
     "170014691C#    ",
     "170014691D#    ",
     "170014691*#    ",
     "170014691#     ",
     "1700146920#    ",
     "1700146921#    ",
     "1700146922#    ",
     "1700146923#    ",
     "1700146924#    ",
     "1700146925#    ",
     "1700146926#    ",
     "1700146927#    ",
     "1700146928#    ",
     "1700146929#    ",
     "170014692A#    ",
     "170014692B#    ",
     "170014692C#    ",
     "170014692D#    ",
     "170014692*#    ",
     "170014692#     ",
     "1700146930#    ",
     "1700146931#    ",
     "1700146932#    ",
     "1700146933#    ",
     "1700146934#    ",
     "1700146935#    ",
     "1700146936#    ",
     "1700146937#    ",
     "1700146938#    ",
     "1700146939#    ",
     "170014693A#    ",
     "170014693B#    ",
     "170014693C#    ",
     "170014693D#    ",
     "170014693*#    ",
     "170014693#     ",
     "1700146940#    ",
     "1700146941#    ",
     "1700146942#    ",
     "1700146943#    ",
     "1700146944#    ",
     "1700146945#    ",
     "1700146946#    ",
     "1700146947#    ",
     "1700146948#    ",
     "1700146949#    ",
     "170014694A#    ",
     "170014694B#    ",
     "170014694C#    ",
     "170014694D#    ",
     "170014694*#    ",
     "170014694#     ",
     "1700146950#    ",
     "1700146951#    ",
     "1700146952#    ",
     "1700146953#    ",
     "1700146954#    ",
     "1700146955#    ",
     "1700146956#    ",
     "1700146957#    ",
     "1700146958#    ",
     "1700146959#    ",
     "170014695A#    ",
     "170014695B#    ",
     "170014695C#    ",
     "170014695D#    ",
     "170014695*#    ",
     "170014695#     ",
     "1700146960#    ",
     "1700146961#    ",
     "1700146962#    ",
     "1700146963#    ",
     "1700146964#    ",
     "1700146965#    ",
     "1700146966#    ",
     "1700146967#    ",
     "1700146968#    ",
     "1700146969#    ",
     "170014696A#    ",
     "170014696B#    ",
     "170014696C#    ",
     "170014696D#    ",
     "170014696*#    ",
     "170014696#     ",
     "1700146970#    ",
     "1700146971#    ",
     "1700146972#    ",
     "1700146973#    ",
     "1700146974#    ",
     "1700146975#    ",
     "1700146976#    ",
     "1700146977#    ",
     "1700146978#    ",
     "1700146979#    ",
     "170014697A#    ",
     "170014697B#    ",
     "170014697C#    ",
     "170014697D#    ",
     "170014697*#    ",
     "170014697#     ",
     "1700146980#    ",
     "1700146981#    ",
     "1700146982#    ",
     "1700146983#    ",
     "1700146984#    ",
     "1700146985#    ",
     "1700146986#    ",
     "1700146987#    ",
     "1700146988#    ",
     "1700146989#    ",
     "170014698A#    ",
     "170014698B#    ",
     "170014698C#    ",
     "170014698D#    ",
     "170014698*#    ",
     "170014698#     ",
     "1700146990#    ",
     "1700146991#    ",
     "1700146992#    ",
     "1700146993#    ",
     "1700146994#    ",
     "1700146995#    ",
     "1700146996#    ",
     "1700146997#    ",
     "1700146998#    ",
     "1700146999#    ",
     "170014699A#    ",
     "170014699B#    ",
     "170014699C#    ",
     "170014699D#    ",
     "170014699*#    ",
     "170014699#     ",
     "17001469A0#    ",
     "17001469A1#    ",
     "17001469A2#    ",
     "17001469A3#    ",
     "17001469A4#    ",
     "17001469A5#    ",
     "17001469A6#    ",
     "17001469A7#    ",
     "17001469A8#    ",
     "17001469A9#    ",
     "17001469AA#    ",
     "17001469AB#    ",
     "17001469AC#    ",
     "17001469AD#    ",
     "17001469A*#    ",
     "17001469A#     ",
     "17001469B0#    ",
     "17001469B1#    ",
     "17001469B2#    ",
     "17001469B3#    ",
     "17001469B4#    ",
     "17001469B5#    ",
     "17001469B6#    ",
     "17001469B7#    ",
     "17001469B8#    ",
     "17001469B9#    ",
     "17001469BA#    ",
     "17001469BB#    ",
     "17001469BC#    ",
     "17001469BD#    ",
     "17001469B*#    ",
     "17001469B#     ",
     "17001469C0#    ",
     "17001469C1#    ",
     "17001469C2#    ",
     "17001469C3#    ",
     "17001469C4#    ",
     "17001469C5#    ",
     "17001469C6#    ",
     "17001469C7#    ",
     "17001469C8#    ",
     "17001469C9#    ",
     "17001469CA#    ",
     "17001469CB#    ",
     "17001469CC#    ",
     "17001469CD#    ",
     "17001469C*#    ",
     "17001469C#     ",
     "17001469D0#    ",
     "17001469D1#    ",
     "17001469D2#    ",
     "17001469D3#    ",
     "17001469D4#    ",
     "17001469D5#    ",
     "17001469D6#    ",
     "17001469D7#    ",
     "17001469D8#    ",
     "17001469D9#    ",
     "17001469DA#    ",
     "17001469DB#    ",
     "17001469DC#    ",
     "17001469DD#    ",
     "17001469D*#    ",
     "17001469D#     ",
     "17001469*0#    ",
     "17001469*1#    ",
     "17001469*2#    ",
     "17001469*3#    ",
     "17001469*4#    ",
     "17001469*5#    ",
     "17001469*6#    ",
     "17001469*7#    ",
     "17001469*8#    ",
     "17001469*9#    ",
     "17001469*A#    ",
     "17001469*B#    ",
     "17001469*C#    ",
     "17001469*D#    ",
     "17001469**#    ",
     "17001469*#     ",
     "01700146915#   ",
     "11700146915#   ",
     "21700146915#   ",
     "31700146915#   ",
     "41700146915#   ",
     "51700146915#   ",
     "61700146915#   ",
     "71700146915#   ",
     "81700146915#   ",
     "91700146915#   ",
     "A1700146915#   ",
     "B1700146915#   ",
     "C1700146915#   ",
     "D1700146915#   ",
     "*1700146915#   ",
     "10700146915#   ",
     "11700146915#   ",
     "12700146915#   ",
     "13700146915#   ",
     "14700146915#   ",
     "15700146915#   ",
     "16700146915#   ",
     "17700146915#   ",
     "18700146915#   ",
     "19700146915#   ",
     "1A700146915#   ",
     "1B700146915#   ",
     "1C700146915#   ",
     "1D700146915#   ",
     "1*700146915#   ",
     "17000146915#   ",
     "17100146915#   ",
     "17200146915#   ",
     "17300146915#   ",
     "17400146915#   ",
     "17500146915#   ",
     "17600146915#   ",
     "17700146915#   ",
     "17800146915#   ",
     "17900146915#   ",
     "17A00146915#   ",
     "17B00146915#   ",
     "17C00146915#   ",
     "17D00146915#   ",
     "17*00146915#   ",
     "17000146915#   ",
     "17010146915#   ",
     "17020146915#   ",
     "17030146915#   ",
     "17040146915#   ",
     "17050146915#   ",
     "17060146915#   ",
     "17070146915#   ",
     "17080146915#   ",
     "17090146915#   ",
     "170A0146915#   ",
     "170B0146915#   ",
     "170C0146915#   ",
     "170D0146915#   ",
     "170*0146915#   ",
     "17000146915#   ",
     "17001146915#   ",
     "17002146915#   ",
     "17003146915#   ",
     "17004146915#   ",
     "17005146915#   ",
     "17006146915#   ",
     "17007146915#   ",
     "17008146915#   ",
     "17009146915#   ",
     "1700A146915#   ",
     "1700B146915#   ",
     "1700C146915#   ",
     "1700D146915#   ",
     "1700*146915#   ",
     "17001046915#   ",
     "17001146915#   ",
     "17001246915#   ",
     "17001346915#   ",
     "17001446915#   ",
     "17001546915#   ",
     "17001646915#   ",
     "17001746915#   ",
     "17001846915#   ",
     "17001946915#   ",
     "17001A46915#   ",
     "17001B46915#   ",
     "17001C46915#   ",
     "17001D46915#   ",
     "17001*46915#   ",
     "17001406915#   ",
     "17001416915#   ",
     "17001426915#   ",
     "17001436915#   ",
     "17001446915#   ",
     "17001456915#   ",
     "17001466915#   ",
     "17001476915#   ",
     "17001486915#   ",
     "17001496915#   ",
     "170014A6915#   ",
     "170014B6915#   ",
     "170014C6915#   ",
     "170014D6915#   ",
     "170014*6915#   ",
     "17001460915#   ",
     "17001461915#   ",
     "17001462915#   ",
     "17001463915#   ",
     "17001464915#   ",
     "17001465915#   ",
     "17001466915#   ",
     "17001467915#   ",
     "17001468915#   ",
     "17001469915#   ",
     "1700146A915#   ",
     "1700146B915#   ",
     "1700146C915#   ",
     "1700146D915#   ",
     "1700146*915#   ",
     "17001469015#   ",
     "17001469115#   ",
     "17001469215#   ",
     "17001469315#   ",
     "17001469415#   ",
     "17001469515#   ",
     "17001469615#   ",
     "17001469715#   ",
     "17001469815#   ",
     "17001469915#   ",
     "17001469A15#   ",
     "17001469B15#   ",
     "17001469C15#   ",
     "17001469D15#   ",
     "17001469*15#   ",
     "17001469105#   ",
     "17001469115#   ",
     "17001469125#   ",
     "17001469135#   ",
     "17001469145#   ",
     "17001469155#   ",
     "17001469165#   ",
     "17001469175#   ",
     "17001469185#   ",
     "17001469195#   ",
     "170014691A5#   ",
     "170014691B5#   ",
     "170014691C5#   ",
     "170014691D5#   ",
     "170014691*5#   ",
     "17001469150#   ",
     "17001469151#   ",
     "17001469152#   ",
     "17001469153#   ",
     "17001469154#   ",
     "17001469155#   ",
     "17001469156#   ",
     "17001469157#   ",
     "17001469158#   ",
     "17001469159#   ",
     "1700146915A#   ",
     "1700146915B#   ",
     "1700146915C#   ",
     "1700146915D#   ",
     "1700146915*#   ",
     "700146915#     ",
     "100146915#     ",
     "170146915#     ",
     "170146915#     ",
     "170046915#     ",
     "170016915#     ",
     "170014915#     ",
     "170014615#     ",
     "170014695#     ",
     "170014691#     ",
     "#              ",
     "1#             ",
     "17#            ",
     "170#           ",
     "1700#          ",
     "17001#         ",
     "170014#        ",
     "1700146#       ",
     "17001469#      ",
     "170014691#     ",
     "1700146915#    ",
     "1700146915#    ",
     "700146915#     ",
     "00146915#      ",
     "0146915#       ",
     "146915#        ",
     "46915#         ",
     "6915#          ",
     "915#           ",
     "15#            ",
     "5#             ",
     "#              ",
     "0550220373#    ",
     "1550220373#    ",
     "2550220373#    ",
     "3550220373#    ",
     "4550220373#    ",
     "5550220373#    ",
     "6550220373#    ",
     "7550220373#    ",
     "8550220373#    ",
     "9550220373#    ",
     "A550220373#    ",
     "B550220373#    ",
     "C550220373#    ",
     "D550220373#    ",
     "*550220373#    ",
     "1050220373#    ",
     "1150220373#    ",
     "1250220373#    ",
     "1350220373#    ",
     "1450220373#    ",
     "1550220373#    ",
     "1650220373#    ",
     "1750220373#    ",
     "1850220373#    ",
     "1950220373#    ",
     "1A50220373#    ",
     "1B50220373#    ",
     "1C50220373#    ",
     "1D50220373#    ",
     "1*50220373#    ",
     "1500220373#    ",
     "1510220373#    ",
     "1520220373#    ",
     "1530220373#    ",
     "1540220373#    ",
     "1550220373#    ",
     "1560220373#    ",
     "1570220373#    ",
     "1580220373#    ",
     "1590220373#    ",
     "15A0220373#    ",
     "15B0220373#    ",
     "15C0220373#    ",
     "15D0220373#    ",
     "15*0220373#    ",
     "1550220373#    ",
     "1551220373#    ",
     "1552220373#    ",
     "1553220373#    ",
     "1554220373#    ",
     "1555220373#    ",
     "1556220373#    ",
     "1557220373#    ",
     "1558220373#    ",
     "1559220373#    ",
     "155A220373#    ",
     "155B220373#    ",
     "155C220373#    ",
     "155D220373#    ",
     "155*220373#    ",
     "1550020373#    ",
     "1550120373#    ",
     "1550220373#    ",
     "1550320373#    ",
     "1550420373#    ",
     "1550520373#    ",
     "1550620373#    ",
     "1550720373#    ",
     "1550820373#    ",
     "1550920373#    ",
     "1550A20373#    ",
     "1550B20373#    ",
     "1550C20373#    ",
     "1550D20373#    ",
     "1550*20373#    ",
     "1550200373#    ",
     "1550210373#    ",
     "1550220373#    ",
     "1550230373#    ",
     "1550240373#    ",
     "1550250373#    ",
     "1550260373#    ",
     "1550270373#    ",
     "1550280373#    ",
     "1550290373#    ",
     "15502A0373#    ",
     "15502B0373#    ",
     "15502C0373#    ",
     "15502D0373#    ",
     "15502*0373#    ",
     "1550220373#    ",
     "1550221373#    ",
     "1550222373#    ",
     "1550223373#    ",
     "1550224373#    ",
     "1550225373#    ",
     "1550226373#    ",
     "1550227373#    ",
     "1550228373#    ",
     "1550229373#    ",
     "155022A373#    ",
     "155022B373#    ",
     "155022C373#    ",
     "155022D373#    ",
     "155022*373#    ",
     "1550220073#    ",
     "1550220173#    ",
     "1550220273#    ",
     "1550220373#    ",
     "1550220473#    ",
     "1550220573#    ",
     "1550220673#    ",
     "1550220773#    ",
     "1550220873#    ",
     "1550220973#    ",
     "1550220A73#    ",
     "1550220B73#    ",
     "1550220C73#    ",
     "1550220D73#    ",
     "1550220*73#    ",
     "1550220303#    ",
     "1550220313#    ",
     "1550220323#    ",
     "1550220333#    ",
     "1550220343#    ",
     "1550220353#    ",
     "1550220363#    ",
     "1550220373#    ",
     "1550220383#    ",
     "1550220393#    ",
     "15502203A3#    ",
     "15502203B3#    ",
     "15502203C3#    ",
     "15502203D3#    ",
     "15502203*3#    ",
     "1550220370#    ",
     "1550220371#    ",
     "1550220372#    ",
     "1550220373#    ",
     "1550220374#    ",
     "1550220375#    ",
     "1550220376#    ",
     "1550220377#    ",
     "1550220378#    ",
     "1550220379#    ",
     "155022037A#    ",
     "155022037B#    ",
     "155022037C#    ",
     "155022037D#    ",
     "155022037*#    ",
     "00#            ",
     "01#            ",
     "02#            ",
     "03#            ",
     "04#            ",
     "05#            ",
     "06#            ",
     "07#            ",
     "08#            ",
     "09#            ",
     "0A#            ",
     "0B#            ",
     "0C#            ",
     "0D#            ",
     "0*#            ",
     "0#             ",
     "10#            ",
     "11#            ",
     "12#            ",
     "13#            ",
     "14#            ",
     "15#            ",
     "16#            ",
     "17#            ",
     "18#            ",
     "19#            ",
     "1A#            ",
     "1B#            ",
     "1C#            ",
     "1D#            ",
     "1*#            ",
     "1#             ",
     "20#            ",
     "21#            ",
     "22#            ",
     "23#            ",
     "24#            ",
     "25#            ",
     "26#            ",
     "27#            ",
     "28#            ",
     "29#            ",
     "2A#            ",
     "2B#            ",
     "2C#            ",
     "2D#            ",
     "2*#            ",
     "2#             ",
     "30#            ",
     "31#            ",
     "32#            ",
     "33#            ",
     "34#            ",
     "35#            ",
     "36#            ",
     "37#            ",
     "38#            ",
     "39#            ",
     "3A#            ",
     "3B#            ",
     "3C#            ",
     "3D#            ",
     "3*#            ",
     "3#             ",
     "40#            ",
     "41#            ",
     "42#            ",
     "43#            ",
     "44#            ",
     "45#            ",
     "46#            ",
     "47#            ",
     "48#            ",
     "49#            ",
     "4A#            ",
     "4B#            ",
     "4C#            ",
     "4D#            ",
     "4*#            ",
     "4#             ",
     "50#            ",
     "51#            ",
     "52#            ",
     "53#            ",
     "54#            ",
     "55#            ",
     "56#            ",
     "57#            ",
     "58#            ",
     "59#            ",
     "5A#            ",
     "5B#            ",
     "5C#            ",
     "5D#            ",
     "5*#            ",
     "5#             ",
     "60#            ",
     "61#            ",
     "62#            ",
     "63#            ",
     "64#            ",
     "65#            ",
     "66#            ",
     "67#            ",
     "68#            ",
     "69#            ",
     "6A#            ",
     "6B#            ",
     "6C#            ",
     "6D#            ",
     "6*#            ",
     "6#             ",
     "70#            ",
     "71#            ",
     "72#            ",
     "73#            ",
     "74#            ",
     "75#            ",
     "76#            ",
     "77#            ",
     "78#            ",
     "79#            ",
     "7A#            ",
     "7B#            ",
     "7C#            ",
     "7D#            ",
     "7*#            ",
     "7#             ",
     "80#            ",
     "81#            ",
     "82#            ",
     "83#            ",
     "84#            ",
     "85#            ",
     "86#            ",
     "87#            ",
     "88#            ",
     "89#            ",
     "8A#            ",
     "8B#            ",
     "8C#            ",
     "8D#            ",
     "8*#            ",
     "8#             ",
     "90#            ",
     "91#            ",
     "92#            ",
     "93#            ",
     "94#            ",
     "95#            ",
     "96#            ",
     "97#            ",
     "98#            ",
     "99#            ",
     "9A#            ",
     "9B#            ",
     "9C#            ",
     "9D#            ",
     "9*#            ",
     "9#             ",
     "A0#            ",
     "A1#            ",
     "A2#            ",
     "A3#            ",
     "A4#            ",
     "A5#            ",
     "A6#            ",
     "A7#            ",
     "A8#            ",
     "A9#            ",
     "AA#            ",
     "AB#            ",
     "AC#            ",
     "AD#            ",
     "A*#            ",
     "A#             ",
     "B0#            ",
     "B1#            ",
     "B2#            ",
     "B3#            ",
     "B4#            ",
     "B5#            ",
     "B6#            ",
     "B7#            ",
     "B8#            ",
     "B9#            ",
     "BA#            ",
     "BB#            ",
     "BC#            ",
     "BD#            ",
     "B*#            ",
     "B#             ",
     "C0#            ",
     "C1#            ",
     "C2#            ",
     "C3#            ",
     "C4#            ",
     "C5#            ",
     "C6#            ",
     "C7#            ",
     "C8#            ",
     "C9#            ",
     "CA#            ",
     "CB#            ",
     "CC#            ",
     "CD#            ",
     "C*#            ",
     "C#             ",
     "D0#            ",
     "D1#            ",
     "D2#            ",
     "D3#            ",
     "D4#            ",
     "D5#            ",
     "D6#            ",
     "D7#            ",
     "D8#            ",
     "D9#            ",
     "DA#            ",
     "DB#            ",
     "DC#            ",
     "DD#            ",
     "D*#            ",
     "D#             ",
     "*0#            ",
     "*1#            ",
     "*2#            ",
     "*3#            ",
     "*4#            ",
     "*5#            ",
     "*6#            ",
     "*7#            ",
     "*8#            ",
     "*9#            ",
     "*A#            ",
     "*B#            ",
     "*C#            ",
     "*D#            ",
     "**#            ",
     "*#             ",
     "1550220300#    ",
     "1550220301#    ",
     "1550220302#    ",
     "1550220303#    ",
     "1550220304#    ",
     "1550220305#    ",
     "1550220306#    ",
     "1550220307#    ",
     "1550220308#    ",
     "1550220309#    ",
     "155022030A#    ",
     "155022030B#    ",
     "155022030C#    ",
     "155022030D#    ",
     "155022030*#    ",
     "155022030#     ",
     "1550220310#    ",
     "1550220311#    ",
     "1550220312#    ",
     "1550220313#    ",
     "1550220314#    ",
     "1550220315#    ",
     "1550220316#    ",
     "1550220317#    ",
     "1550220318#    ",
     "1550220319#    ",
     "155022031A#    ",
     "155022031B#    ",
     "155022031C#    ",
     "155022031D#    ",
     "155022031*#    ",
     "155022031#     ",
     "1550220320#    ",
     "1550220321#    ",
     "1550220322#    ",
     "1550220323#    ",
     "1550220324#    ",
     "1550220325#    ",
     "1550220326#    ",
     "1550220327#    ",
     "1550220328#    ",
     "1550220329#    ",
     "155022032A#    ",
     "155022032B#    ",
     "155022032C#    ",
     "155022032D#    ",
     "155022032*#    ",
     "155022032#     ",
     "1550220330#    ",
     "1550220331#    ",
     "1550220332#    ",
     "1550220333#    ",
     "1550220334#    ",
     "1550220335#    ",
     "1550220336#    ",
     "1550220337#    ",
     "1550220338#    ",
     "1550220339#    ",
     "155022033A#    ",
     "155022033B#    ",
     "155022033C#    ",
     "155022033D#    ",
     "155022033*#    ",
     "155022033#     ",
     "1550220340#    ",
     "1550220341#    ",
     "1550220342#    ",
     "1550220343#    ",
     "1550220344#    ",
     "1550220345#    ",
     "1550220346#    ",
     "1550220347#    ",
     "1550220348#    ",
     "1550220349#    ",
     "155022034A#    ",
     "155022034B#    ",
     "155022034C#    ",
     "155022034D#    ",
     "155022034*#    ",
     "155022034#     ",
     "1550220350#    ",
     "1550220351#    ",
     "1550220352#    ",
     "1550220353#    ",
     "1550220354#    ",
     "1550220355#    ",
     "1550220356#    ",
     "1550220357#    ",
     "1550220358#    ",
     "1550220359#    ",
     "155022035A#    ",
     "155022035B#    ",
     "155022035C#    ",
     "155022035D#    ",
     "155022035*#    ",
     "155022035#     ",
     "1550220360#    ",
     "1550220361#    ",
     "1550220362#    ",
     "1550220363#    ",
     "1550220364#    ",
     "1550220365#    ",
     "1550220366#    ",
     "1550220367#    ",
     "1550220368#    ",
     "1550220369#    ",
     "155022036A#    ",
     "155022036B#    ",
     "155022036C#    ",
     "155022036D#    ",
     "155022036*#    ",
     "155022036#     ",
     "1550220370#    ",
     "1550220371#    ",
     "1550220372#    ",
     "1550220373#    ",
     "1550220374#    ",
     "1550220375#    ",
     "1550220376#    ",
     "1550220377#    ",
     "1550220378#    ",
     "1550220379#    ",
     "155022037A#    ",
     "155022037B#    ",
     "155022037C#    ",
     "155022037D#    ",
     "155022037*#    ",
     "155022037#     ",
     "1550220380#    ",
     "1550220381#    ",
     "1550220382#    ",
     "1550220383#    ",
     "1550220384#    ",
     "1550220385#    ",
     "1550220386#    ",
     "1550220387#    ",
     "1550220388#    ",
     "1550220389#    ",
     "155022038A#    ",
     "155022038B#    ",
     "155022038C#    ",
     "155022038D#    ",
     "155022038*#    ",
     "155022038#     ",
     "1550220390#    ",
     "1550220391#    ",
     "1550220392#    ",
     "1550220393#    ",
     "1550220394#    ",
     "1550220395#    ",
     "1550220396#    ",
     "1550220397#    ",
     "1550220398#    ",
     "1550220399#    ",
     "155022039A#    ",
     "155022039B#    ",
     "155022039C#    ",
     "155022039D#    ",
     "155022039*#    ",
     "155022039#     ",
     "15502203A0#    ",
     "15502203A1#    ",
     "15502203A2#    ",
     "15502203A3#    ",
     "15502203A4#    ",
     "15502203A5#    ",
     "15502203A6#    ",
     "15502203A7#    ",
     "15502203A8#    ",
     "15502203A9#    ",
     "15502203AA#    ",
     "15502203AB#    ",
     "15502203AC#    ",
     "15502203AD#    ",
     "15502203A*#    ",
     "15502203A#     ",
     "15502203B0#    ",
     "15502203B1#    ",
     "15502203B2#    ",
     "15502203B3#    ",
     "15502203B4#    ",
     "15502203B5#    ",
     "15502203B6#    ",
     "15502203B7#    ",
     "15502203B8#    ",
     "15502203B9#    ",
     "15502203BA#    ",
     "15502203BB#    ",
     "15502203BC#    ",
     "15502203BD#    ",
     "15502203B*#    ",
     "15502203B#     ",
     "15502203C0#    ",
     "15502203C1#    ",
     "15502203C2#    ",
     "15502203C3#    ",
     "15502203C4#    ",
     "15502203C5#    ",
     "15502203C6#    ",
     "15502203C7#    ",
     "15502203C8#    ",
     "15502203C9#    ",
     "15502203CA#    ",
     "15502203CB#    ",
     "15502203CC#    ",
     "15502203CD#    ",
     "15502203C*#    ",
     "15502203C#     ",
     "15502203D0#    ",
     "15502203D1#    ",
     "15502203D2#    ",
     "15502203D3#    ",
     "15502203D4#    ",
     "15502203D5#    ",
     "15502203D6#    ",
     "15502203D7#    ",
     "15502203D8#    ",
     "15502203D9#    ",
     "15502203DA#    ",
     "15502203DB#    ",
     "15502203DC#    ",
     "15502203DD#    ",
     "15502203D*#    ",
     "15502203D#     ",
     "15502203*0#    ",
     "15502203*1#    ",
     "15502203*2#    ",
     "15502203*3#    ",
     "15502203*4#    ",
     "15502203*5#    ",
     "15502203*6#    ",
     "15502203*7#    ",
     "15502203*8#    ",
     "15502203*9#    ",
     "15502203*A#    ",
     "15502203*B#    ",
     "15502203*C#    ",
     "15502203*D#    ",
     "15502203**#    ",
     "15502203*#     ",
     "01550220373#   ",
     "11550220373#   ",
     "21550220373#   ",
     "31550220373#   ",
     "41550220373#   ",
     "51550220373#   ",
     "61550220373#   ",
     "71550220373#   ",
     "81550220373#   ",
     "91550220373#   ",
     "A1550220373#   ",
     "B1550220373#   ",
     "C1550220373#   ",
     "D1550220373#   ",
     "*1550220373#   ",
     "10550220373#   ",
     "11550220373#   ",
     "12550220373#   ",
     "13550220373#   ",
     "14550220373#   ",
     "15550220373#   ",
     "16550220373#   ",
     "17550220373#   ",
     "18550220373#   ",
     "19550220373#   ",
     "1A550220373#   ",
     "1B550220373#   ",
     "1C550220373#   ",
     "1D550220373#   ",
     "1*550220373#   ",
     "15050220373#   ",
     "15150220373#   ",
     "15250220373#   ",
     "15350220373#   ",
     "15450220373#   ",
     "15550220373#   ",
     "15650220373#   ",
     "15750220373#   ",
     "15850220373#   ",
     "15950220373#   ",
     "15A50220373#   ",
     "15B50220373#   ",
     "15C50220373#   ",
     "15D50220373#   ",
     "15*50220373#   ",
     "15500220373#   ",
     "15510220373#   ",
     "15520220373#   ",
     "15530220373#   ",
     "15540220373#   ",
     "15550220373#   ",
     "15560220373#   ",
     "15570220373#   ",
     "15580220373#   ",
     "15590220373#   ",
     "155A0220373#   ",
     "155B0220373#   ",
     "155C0220373#   ",
     "155D0220373#   ",
     "155*0220373#   ",
     "15500220373#   ",
     "15501220373#   ",
     "15502220373#   ",
     "15503220373#   ",
     "15504220373#   ",
     "15505220373#   ",
     "15506220373#   ",
     "15507220373#   ",
     "15508220373#   ",
     "15509220373#   ",
     "1550A220373#   ",
     "1550B220373#   ",
     "1550C220373#   ",
     "1550D220373#   ",
     "1550*220373#   ",
     "15502020373#   ",
     "15502120373#   ",
     "15502220373#   ",
     "15502320373#   ",
     "15502420373#   ",
     "15502520373#   ",
     "15502620373#   ",
     "15502720373#   ",
     "15502820373#   ",
     "15502920373#   ",
     "15502A20373#   ",
     "15502B20373#   ",
     "15502C20373#   ",
     "15502D20373#   ",
     "15502*20373#   ",
     "15502200373#   ",
     "15502210373#   ",
     "15502220373#   ",
     "15502230373#   ",
     "15502240373#   ",
     "15502250373#   ",
     "15502260373#   ",
     "15502270373#   ",
     "15502280373#   ",
     "15502290373#   ",
     "155022A0373#   ",
     "155022B0373#   ",
     "155022C0373#   ",
     "155022D0373#   ",
     "155022*0373#   ",
     "15502200373#   ",
     "15502201373#   ",
     "15502202373#   ",
     "15502203373#   ",
     "15502204373#   ",
     "15502205373#   ",
     "15502206373#   ",
     "15502207373#   ",
     "15502208373#   ",
     "15502209373#   ",
     "1550220A373#   ",
     "1550220B373#   ",
     "1550220C373#   ",
     "1550220D373#   ",
     "1550220*373#   ",
     "15502203073#   ",
     "15502203173#   ",
     "15502203273#   ",
     "15502203373#   ",
     "15502203473#   ",
     "15502203573#   ",
     "15502203673#   ",
     "15502203773#   ",
     "15502203873#   ",
     "15502203973#   ",
     "15502203A73#   ",
     "15502203B73#   ",
     "15502203C73#   ",
     "15502203D73#   ",
     "15502203*73#   ",
     "15502203703#   ",
     "15502203713#   ",
     "15502203723#   ",
     "15502203733#   ",
     "15502203743#   ",
     "15502203753#   ",
     "15502203763#   ",
     "15502203773#   ",
     "15502203783#   ",
     "15502203793#   ",
     "155022037A3#   ",
     "155022037B3#   ",
     "155022037C3#   ",
     "155022037D3#   ",
     "155022037*3#   ",
     "15502203730#   ",
     "15502203731#   ",
     "15502203732#   ",
     "15502203733#   ",
     "15502203734#   ",
     "15502203735#   ",
     "15502203736#   ",
     "15502203737#   ",
     "15502203738#   ",
     "15502203739#   ",
     "1550220373A#   ",
     "1550220373B#   ",
     "1550220373C#   ",
     "1550220373D#   ",
     "1550220373*#   ",
     "550220373#     ",
     "150220373#     ",
     "150220373#     ",
     "155220373#     ",
     "155020373#     ",
     "155020373#     ",
     "155022373#     ",
     "155022073#     ",
     "155022033#     ",
     "155022037#     ",
     "#              ",
     "1#             ",
     "15#            ",
     "155#           ",
     "1550#          ",
     "15502#         ",
     "155022#        ",
     "1550220#       ",
     "15502203#      ",
     "155022037#     ",
     "1550220373#    ",
     "1550220373#    ",
     "550220373#     ",
     "50220373#      ",
     "0220373#       ",
     "220373#        ",
     "20373#         ",
     "0373#          ",
     "373#           ",
     "73#            ",
     "3#             ",
     "#              ",
     "1700146915#    ",
     "1700146915#    ",
     "1500146915#    ",
     "1550146915#    ",
     "1550146915#    ",
     "1550246915#    ",
     "1550226915#    ",
     "1550220915#    ",
     "1550220315#    ",
     "1550220375#    ",
     "1550220373#    ",
     "1550220373#    ",
     "1550220373#    ",
     "1750220373#    ",
     "1700220373#    ",
     "1700220373#    ",
     "1700120373#    ",
     "1700140373#    ",
     "1700146373#    ",
     "1700146973#    ",
     "1700146913#    ",
     "1700146915#    "
   ); 

end testbench_pkg;

package body testbench_pkg is
end testbench_pkg;
