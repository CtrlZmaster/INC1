library IEEE;
use IEEE.std_logic_1164.all;

package testbench_pkg is
   constant FILE_NAME : string := "chk_sim_sig_basic.txt";

   constant N_TEST_WORDS : integer := 48; 
   type t_test_words     is array (1 to N_TEST_WORDS) 
                                  of string(1 to 15);
   constant test_words : t_test_words :=
   ( 
     "1700146915#    ",
     "1234567890*#   ",
     "1700146915#    ",
     "234567890*#    ",
     "1700146915#    ",
     "34567890*#     ",
     "1700146915#    ",
     "4567890*#      ",
     "1700146915#    ",
     "567890*#       ",
     "1700146915#    ",
     "67890*#        ",
     "1700146915#    ",
     "7890*#         ",
     "1700146915#    ",
     "890*#          ",
     "1700146915#    ",
     "90*#           ",
     "1700146915#    ",
     "0*#            ",
     "1700146915#    ",
     "*#             ",
     "1700146915#    ",
     "#              ",
     "1550220373#    ",
     "1234567890*#   ",
     "1550220373#    ",
     "234567890*#    ",
     "1550220373#    ",
     "34567890*#     ",
     "1550220373#    ",
     "4567890*#      ",
     "1550220373#    ",
     "567890*#       ",
     "1550220373#    ",
     "67890*#        ",
     "1550220373#    ",
     "7890*#         ",
     "1550220373#    ",
     "890*#          ",
     "1550220373#    ",
     "90*#           ",
     "1550220373#    ",
     "0*#            ",
     "1550220373#    ",
     "*#             ",
     "1550220373#    ",
     "#              "
   ); 

end testbench_pkg;

package body testbench_pkg is
end testbench_pkg;
